module top ( a , c ); wire a ; wire c;
    input a;
    output c;
 
    assign c = a;

endmodule
